----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Reed Foster
-- 
-- Create Date:    21:55:39 04/07/2016 
-- Design Name: 
-- Module Name:    rom64x8 - behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
-- 64B read only memory
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom4kB is
   port (addr     : in  std_logic_vector (11 downto 0);
         sel      : in  std_logic;
         data_out : out std_logic_vector (7 downto 0);
         out_ctl  : out std_logic
	);
end rom4kB;

architecture behavioral of rom4kB is
   type array_type is array (0 to 4095) of std_logic_vector (7 downto 0);
   type prog_type is array (0 to 1023) of std_logic_vector (15 downto 0);
   type data_type is array (0 to 2047) of std_logic_vector (7 downto 0);
   constant prog_instr : prog_type := (
--	   fill with desired program (max 1023 instructions)
----------------------------------------------------------------------------------------------------------
--		current program : draw a buffer to ssd1306 oled controller (commented code sends commands to processor)
      0 => x"7eff",
      1 => x"5601",
      2 => x"81ff",
      3 => x"0a27",
      4 => x"c1ff",
      5 => x"56fe",
      6 => x"81ff",
      7 => x"0a26",
      8 => x"c1ff",
      9 => x"660a",
      10 => x"5e01",
      11 => x"4e00",
      12 => x"2143",
      13 => x"5006",
      14 => x"0b22",
      15 => x"40f8",
      16 => x"0000",
      17 => x"5601",
      18 => x"81ff",
      19 => x"0a27",
      20 => x"c1ff",
      21 => x"56e7",
      22 => x"81ff",
      23 => x"0a26",
      24 => x"c1ff",
      25 => x"567f",
      26 => x"81ff",
      27 => x"0a26",
      28 => x"c1ff",
      29 => x"661f",
      30 => x"5e01",
      31 => x"4e00",
      32 => x"2143",
      33 => x"502a",
      34 => x"7e0c",
      35 => x"8d00",
      36 => x"7eff",
      37 => x"c5fe",
      38 => x"7604",
      39 => x"85ff",
      40 => x"2ea7",
      41 => x"c5ff",
      42 => x"7640",
      43 => x"85ff",
      44 => x"2ea6",
      45 => x"6906",
      46 => x"0000",
      47 => x"40f6",
      48 => x"0000",
      49 => x"76fb",
      50 => x"85ff",
      51 => x"2ea6",
      52 => x"c5ff",
      53 => x"40d4",
      54 => x"0b22",
      55 => x"7eff",
      56 => x"7620",
      57 => x"85ff",
      58 => x"2ea6",
      59 => x"6906",
      60 => x"0000",
      61 => x"40f6",
      62 => x"0000",
      63 => x"5680",
      64 => x"81ff",
      65 => x"0a27",
      66 => x"c1ff",
      67 => x"7e08",
      68 => x"5e01",
      69 => x"4e08",
      70 => x"660c",
      71 => x"21a3",
      72 => x"683a",
      73 => x"0000",
      74 => x"66ff",
      75 => x"5600",
      76 => x"22a3",
      77 => x"682c",
      78 => x"0000",
      79 => x"9500",
      80 => x"7eff",
      81 => x"c5fe",
      82 => x"7604",
      83 => x"85ff",
      84 => x"2ea7",
      85 => x"c5ff",
      86 => x"7640",
      87 => x"85ff",
      88 => x"2ea6",
      89 => x"6906",
      90 => x"0000",
      91 => x"40f6",
      92 => x"0000",
      93 => x"76fb",
      94 => x"85ff",
      95 => x"2ea6",
      96 => x"c5ff",
      97 => x"08e2",
      98 => x"40d2",
      99 => x"1342",
      100 => x"40c2",
      101 => x"0b22",
      102 => x"0000",
      103 => x"40fe",
      others => x"0000"

   );
   constant prog_data : data_type := (
      --fill with data to be used in program
      --data
      0    => x"00", 1    => x"00", 2    => x"00", 3    => x"00", 4    => x"00", 5    => x"00", 6    => x"00", 7    => x"00", 8    => x"00", 9    => x"00", 10   => x"00", 11   => x"00", 12   => x"00", 13   => x"00", 14   => x"00", 15   => x"00",
      16   => x"00", 17   => x"00", 18   => x"00", 19   => x"00", 20   => x"00", 21   => x"00", 22   => x"00", 23   => x"00", 24   => x"00", 25   => x"00", 26   => x"00", 27   => x"00", 28   => x"00", 29   => x"00", 30   => x"00", 31   => x"00",
      32   => x"00", 33   => x"00", 34   => x"00", 35   => x"00", 36   => x"00", 37   => x"00", 38   => x"00", 39   => x"00", 40   => x"00", 41   => x"00", 42   => x"00", 43   => x"00", 44   => x"00", 45   => x"00", 46   => x"00", 47   => x"00",
      48   => x"00", 49   => x"00", 50   => x"00", 51   => x"00", 52   => x"00", 53   => x"00", 54   => x"00", 55   => x"00", 56   => x"00", 57   => x"00", 58   => x"00", 59   => x"00", 60   => x"00", 61   => x"00", 62   => x"00", 63   => x"00",
      64   => x"00", 65   => x"00", 66   => x"00", 67   => x"00", 68   => x"00", 69   => x"00", 70   => x"00", 71   => x"00", 72   => x"00", 73   => x"00", 74   => x"00", 75   => x"00", 76   => x"00", 77   => x"00", 78   => x"00", 79   => x"00",
      80   => x"00", 81   => x"00", 82   => x"00", 83   => x"00", 84   => x"00", 85   => x"00", 86   => x"00", 87   => x"00", 88   => x"00", 89   => x"00", 90   => x"00", 91   => x"00", 92   => x"00", 93   => x"00", 94   => x"00", 95   => x"00",
      96   => x"00", 97   => x"00", 98   => x"00", 99   => x"00", 100  => x"00", 101  => x"00", 102  => x"00", 103  => x"00", 104  => x"00", 105  => x"00", 106  => x"00", 107  => x"00", 108  => x"00", 109  => x"00", 110  => x"00", 111  => x"00",
      112  => x"00", 113  => x"00", 114  => x"00", 115  => x"00", 116  => x"00", 117  => x"00", 118  => x"00", 119  => x"00", 120  => x"00", 121  => x"00", 122  => x"00", 123  => x"00", 124  => x"00", 125  => x"00", 126  => x"00", 127  => x"00",
      128  => x"00", 129  => x"00", 130  => x"00", 131  => x"00", 132  => x"00", 133  => x"00", 134  => x"00", 135  => x"00", 136  => x"00", 137  => x"00", 138  => x"00", 139  => x"00", 140  => x"00", 141  => x"00", 142  => x"00", 143  => x"00",
      144  => x"00", 145  => x"00", 146  => x"00", 147  => x"00", 148  => x"00", 149  => x"00", 150  => x"00", 151  => x"00", 152  => x"00", 153  => x"00", 154  => x"00", 155  => x"00", 156  => x"00", 157  => x"00", 158  => x"00", 159  => x"00",
      160  => x"00", 161  => x"00", 162  => x"00", 163  => x"00", 164  => x"00", 165  => x"00", 166  => x"00", 167  => x"00", 168  => x"00", 169  => x"00", 170  => x"00", 171  => x"00", 172  => x"00", 173  => x"00", 174  => x"00", 175  => x"00",
      176  => x"00", 177  => x"00", 178  => x"00", 179  => x"00", 180  => x"00", 181  => x"00", 182  => x"00", 183  => x"00", 184  => x"00", 185  => x"00", 186  => x"00", 187  => x"00", 188  => x"00", 189  => x"00", 190  => x"00", 191  => x"00",
      192  => x"00", 193  => x"00", 194  => x"00", 195  => x"00", 196  => x"00", 197  => x"00", 198  => x"00", 199  => x"00", 200  => x"00", 201  => x"00", 202  => x"00", 203  => x"00", 204  => x"00", 205  => x"00", 206  => x"00", 207  => x"00",
      208  => x"00", 209  => x"00", 210  => x"00", 211  => x"00", 212  => x"00", 213  => x"00", 214  => x"00", 215  => x"00", 216  => x"00", 217  => x"00", 218  => x"00", 219  => x"00", 220  => x"00", 221  => x"00", 222  => x"00", 223  => x"00",
      224  => x"00", 225  => x"00", 226  => x"00", 227  => x"00", 228  => x"00", 229  => x"00", 230  => x"00", 231  => x"00", 232  => x"00", 233  => x"00", 234  => x"00", 235  => x"03", 236  => x"00", 237  => x"03", 238  => x"00", 239  => x"00",
      240  => x"30", 241  => x"30", 242  => x"00", 243  => x"00", 244  => x"00", 245  => x"00", 246  => x"00", 247  => x"fc", 248  => x"63", 249  => x"00", 250  => x"00", 251  => x"03", 252  => x"00", 253  => x"03", 254  => x"00", 255  => x"00",
      256  => x"30", 257  => x"30", 258  => x"00", 259  => x"00", 260  => x"00", 261  => x"00", 262  => x"00", 263  => x"fc", 264  => x"67", 265  => x"00", 266  => x"0c", 267  => x"03", 268  => x"00", 269  => x"03", 270  => x"00", 271  => x"00",
      272  => x"30", 273  => x"30", 274  => x"00", 275  => x"00", 276  => x"00", 277  => x"00", 278  => x"00", 279  => x"0c", 280  => x"06", 281  => x"00", 282  => x"0c", 283  => x"03", 284  => x"00", 285  => x"03", 286  => x"00", 287  => x"00",
      288  => x"30", 289  => x"30", 290  => x"3e", 291  => x"76", 292  => x"d8", 293  => x"31", 294  => x"18", 295  => x"0c", 296  => x"66", 297  => x"6c", 298  => x"3e", 299  => x"7b", 300  => x"70", 301  => x"e3", 302  => x"33", 303  => x"18",
      304  => x"30", 305  => x"30", 306  => x"7f", 307  => x"fe", 308  => x"f8", 309  => x"33", 310  => x"18", 311  => x"0c", 312  => x"66", 313  => x"7c", 314  => x"3e", 315  => x"ff", 316  => x"f8", 317  => x"f3", 318  => x"37", 319  => x"18",
      320  => x"f0", 321  => x"3f", 322  => x"61", 323  => x"ce", 324  => x"39", 325  => x"67", 326  => x"0c", 327  => x"fc", 328  => x"63", 329  => x"1c", 330  => x"0c", 331  => x"c7", 332  => x"9c", 333  => x"13", 334  => x"66", 335  => x"0c",
      336  => x"f0", 337  => x"3f", 338  => x"60", 339  => x"86", 340  => x"19", 341  => x"66", 342  => x"0c", 343  => x"fc", 344  => x"67", 345  => x"0c", 346  => x"0c", 347  => x"c3", 348  => x"0c", 349  => x"03", 350  => x"66", 351  => x"0c",
      352  => x"30", 353  => x"30", 354  => x"7e", 355  => x"86", 356  => x"19", 357  => x"66", 358  => x"0c", 359  => x"0c", 360  => x"66", 361  => x"0c", 362  => x"0c", 363  => x"c3", 364  => x"0c", 365  => x"e3", 366  => x"67", 367  => x"0c",
      368  => x"30", 369  => x"30", 370  => x"63", 371  => x"86", 372  => x"19", 373  => x"c6", 374  => x"06", 375  => x"0c", 376  => x"66", 377  => x"0c", 378  => x"0c", 379  => x"c3", 380  => x"0c", 381  => x"33", 382  => x"c6", 383  => x"06",
      384  => x"30", 385  => x"30", 386  => x"63", 387  => x"ce", 388  => x"39", 389  => x"c7", 390  => x"06", 391  => x"0c", 392  => x"66", 393  => x"0c", 394  => x"0c", 395  => x"c3", 396  => x"9c", 397  => x"33", 398  => x"c6", 399  => x"06",
      400  => x"30", 401  => x"30", 402  => x"7f", 403  => x"fe", 404  => x"f8", 405  => x"83", 406  => x"03", 407  => x"fc", 408  => x"67", 409  => x"0c", 410  => x"3c", 411  => x"c3", 412  => x"f8", 413  => x"f3", 414  => x"87", 415  => x"03",
      416  => x"30", 417  => x"30", 418  => x"6e", 419  => x"76", 420  => x"d8", 421  => x"01", 422  => x"03", 423  => x"fc", 424  => x"63", 425  => x"0c", 426  => x"38", 427  => x"c3", 428  => x"70", 429  => x"e3", 430  => x"06", 431  => x"03",
      432  => x"00", 433  => x"00", 434  => x"00", 435  => x"06", 436  => x"18", 437  => x"00", 438  => x"03", 439  => x"00", 440  => x"00", 441  => x"00", 442  => x"00", 443  => x"00", 444  => x"00", 445  => x"00", 446  => x"00", 447  => x"03",
      448  => x"00", 449  => x"00", 450  => x"00", 451  => x"06", 452  => x"18", 453  => x"80", 454  => x"01", 455  => x"00", 456  => x"00", 457  => x"00", 458  => x"00", 459  => x"00", 460  => x"00", 461  => x"00", 462  => x"80", 463  => x"01",
      464  => x"00", 465  => x"00", 466  => x"00", 467  => x"06", 468  => x"18", 469  => x"80", 470  => x"01", 471  => x"00", 472  => x"00", 473  => x"00", 474  => x"00", 475  => x"00", 476  => x"00", 477  => x"00", 478  => x"80", 479  => x"01",
      480  => x"00", 481  => x"00", 482  => x"00", 483  => x"00", 484  => x"00", 485  => x"00", 486  => x"00", 487  => x"00", 488  => x"00", 489  => x"00", 490  => x"00", 491  => x"00", 492  => x"00", 493  => x"00", 494  => x"00", 495  => x"00",
      496  => x"00", 497  => x"00", 498  => x"00", 499  => x"00", 500  => x"00", 501  => x"00", 502  => x"00", 503  => x"00", 504  => x"00", 505  => x"00", 506  => x"00", 507  => x"00", 508  => x"00", 509  => x"00", 510  => x"00", 511  => x"00",
      512  => x"00", 513  => x"00", 514  => x"00", 515  => x"00", 516  => x"00", 517  => x"00", 518  => x"00", 519  => x"00", 520  => x"00", 521  => x"00", 522  => x"00", 523  => x"00", 524  => x"00", 525  => x"00", 526  => x"00", 527  => x"00",
      528  => x"00", 529  => x"00", 530  => x"00", 531  => x"00", 532  => x"00", 533  => x"00", 534  => x"00", 535  => x"00", 536  => x"00", 537  => x"00", 538  => x"00", 539  => x"00", 540  => x"00", 541  => x"00", 542  => x"00", 543  => x"00",
      544  => x"00", 545  => x"00", 546  => x"00", 547  => x"00", 548  => x"00", 549  => x"00", 550  => x"00", 551  => x"00", 552  => x"00", 553  => x"c6", 554  => x"00", 555  => x"00", 556  => x"00", 557  => x"00", 558  => x"00", 559  => x"00",
      560  => x"00", 561  => x"00", 562  => x"00", 563  => x"00", 564  => x"00", 565  => x"c0", 566  => x"1f", 567  => x"00", 568  => x"00", 569  => x"c6", 570  => x"00", 571  => x"00", 572  => x"00", 573  => x"00", 574  => x"00", 575  => x"00",
      576  => x"00", 577  => x"00", 578  => x"00", 579  => x"00", 580  => x"00", 581  => x"c0", 582  => x"7f", 583  => x"00", 584  => x"00", 585  => x"c6", 586  => x"00", 587  => x"00", 588  => x"00", 589  => x"00", 590  => x"00", 591  => x"00",
      592  => x"00", 593  => x"00", 594  => x"00", 595  => x"00", 596  => x"00", 597  => x"c0", 598  => x"60", 599  => x"00", 600  => x"00", 601  => x"c6", 602  => x"00", 603  => x"00", 604  => x"00", 605  => x"00", 606  => x"00", 607  => x"00",
      608  => x"00", 609  => x"00", 610  => x"00", 611  => x"00", 612  => x"00", 613  => x"c0", 614  => x"c0", 615  => x"f8", 616  => x"e0", 617  => x"c6", 618  => x"00", 619  => x"00", 620  => x"00", 621  => x"00", 622  => x"00", 623  => x"00",
      624  => x"00", 625  => x"00", 626  => x"00", 627  => x"00", 628  => x"00", 629  => x"c0", 630  => x"c0", 631  => x"fc", 632  => x"f1", 633  => x"c7", 634  => x"00", 635  => x"00", 636  => x"00", 637  => x"00", 638  => x"00", 639  => x"00",
      640  => x"00", 641  => x"00", 642  => x"00", 643  => x"00", 644  => x"00", 645  => x"c0", 646  => x"c0", 647  => x"84", 648  => x"39", 649  => x"c7", 650  => x"00", 651  => x"00", 652  => x"00", 653  => x"00", 654  => x"00", 655  => x"00",
      656  => x"00", 657  => x"00", 658  => x"00", 659  => x"00", 660  => x"00", 661  => x"c0", 662  => x"c0", 663  => x"80", 664  => x"19", 665  => x"c6", 666  => x"00", 667  => x"00", 668  => x"00", 669  => x"00", 670  => x"00", 671  => x"00",
      672  => x"00", 673  => x"00", 674  => x"00", 675  => x"00", 676  => x"00", 677  => x"c0", 678  => x"c0", 679  => x"f8", 680  => x"19", 681  => x"c6", 682  => x"00", 683  => x"00", 684  => x"00", 685  => x"00", 686  => x"00", 687  => x"00",
      688  => x"00", 689  => x"00", 690  => x"00", 691  => x"00", 692  => x"00", 693  => x"c0", 694  => x"c0", 695  => x"8c", 696  => x"19", 697  => x"c6", 698  => x"00", 699  => x"00", 700  => x"00", 701  => x"00", 702  => x"00", 703  => x"00",
      704  => x"00", 705  => x"00", 706  => x"00", 707  => x"00", 708  => x"00", 709  => x"c0", 710  => x"60", 711  => x"8c", 712  => x"39", 713  => x"07", 714  => x"00", 715  => x"00", 716  => x"00", 717  => x"00", 718  => x"00", 719  => x"00",
      720  => x"00", 721  => x"00", 722  => x"00", 723  => x"00", 724  => x"00", 725  => x"c0", 726  => x"7f", 727  => x"fc", 728  => x"f1", 729  => x"c7", 730  => x"00", 731  => x"00", 732  => x"00", 733  => x"00", 734  => x"00", 735  => x"00",
      736  => x"00", 737  => x"00", 738  => x"00", 739  => x"00", 740  => x"00", 741  => x"c0", 742  => x"1f", 743  => x"b8", 744  => x"e1", 745  => x"c6", 746  => x"00", 747  => x"00", 748  => x"00", 749  => x"00", 750  => x"00", 751  => x"00",
      752  => x"00", 753  => x"00", 754  => x"00", 755  => x"00", 756  => x"00", 757  => x"00", 758  => x"00", 759  => x"00", 760  => x"00", 761  => x"00", 762  => x"00", 763  => x"00", 764  => x"00", 765  => x"00", 766  => x"00", 767  => x"00",
      768  => x"00", 769  => x"00", 770  => x"00", 771  => x"00", 772  => x"00", 773  => x"00", 774  => x"00", 775  => x"00", 776  => x"00", 777  => x"00", 778  => x"00", 779  => x"00", 780  => x"00", 781  => x"00", 782  => x"00", 783  => x"00",
      784  => x"00", 785  => x"00", 786  => x"00", 787  => x"00", 788  => x"00", 789  => x"00", 790  => x"00", 791  => x"00", 792  => x"00", 793  => x"00", 794  => x"00", 795  => x"00", 796  => x"00", 797  => x"00", 798  => x"00", 799  => x"00",
      800  => x"00", 801  => x"00", 802  => x"00", 803  => x"00", 804  => x"00", 805  => x"00", 806  => x"00", 807  => x"00", 808  => x"00", 809  => x"00", 810  => x"00", 811  => x"00", 812  => x"00", 813  => x"00", 814  => x"00", 815  => x"00",
      816  => x"00", 817  => x"00", 818  => x"00", 819  => x"00", 820  => x"00", 821  => x"00", 822  => x"00", 823  => x"00", 824  => x"00", 825  => x"00", 826  => x"00", 827  => x"00", 828  => x"00", 829  => x"00", 830  => x"00", 831  => x"00",
      832  => x"00", 833  => x"00", 834  => x"00", 835  => x"00", 836  => x"00", 837  => x"00", 838  => x"60", 839  => x"80", 840  => x"01", 841  => x"00", 842  => x"00", 843  => x"d8", 844  => x"27", 845  => x"02", 846  => x"00", 847  => x"00",
      848  => x"00", 849  => x"00", 850  => x"00", 851  => x"00", 852  => x"00", 853  => x"00", 854  => x"40", 855  => x"00", 856  => x"01", 857  => x"00", 858  => x"00", 859  => x"64", 860  => x"29", 861  => x"02", 862  => x"00", 863  => x"00",
      864  => x"00", 865  => x"00", 866  => x"00", 867  => x"00", 868  => x"00", 869  => x"02", 870  => x"40", 871  => x"00", 872  => x"01", 873  => x"00", 874  => x"44", 875  => x"42", 876  => x"29", 877  => x"02", 878  => x"00", 879  => x"00",
      880  => x"f0", 881  => x"98", 882  => x"86", 883  => x"d1", 884  => x"0c", 885  => x"87", 886  => x"71", 887  => x"00", 888  => x"67", 889  => x"03", 890  => x"44", 891  => x"02", 892  => x"29", 893  => x"02", 894  => x"00", 895  => x"00",
      896  => x"48", 897  => x"24", 898  => x"49", 899  => x"22", 900  => x"12", 901  => x"42", 902  => x"4a", 903  => x"00", 904  => x"49", 905  => x"01", 906  => x"44", 907  => x"02", 908  => x"27", 909  => x"02", 910  => x"00", 911  => x"00",
      912  => x"30", 913  => x"3c", 914  => x"c9", 915  => x"23", 916  => x"1c", 917  => x"c2", 918  => x"4b", 919  => x"00", 920  => x"49", 921  => x"01", 922  => x"44", 923  => x"02", 924  => x"21", 925  => x"02", 926  => x"00", 927  => x"00",
      928  => x"08", 929  => x"04", 930  => x"49", 931  => x"20", 932  => x"12", 933  => x"42", 934  => x"48", 935  => x"00", 936  => x"89", 937  => x"01", 938  => x"44", 939  => x"44", 940  => x"21", 941  => x"02", 942  => x"00", 943  => x"00",
      944  => x"78", 945  => x"38", 946  => x"89", 947  => x"73", 948  => x"3c", 949  => x"84", 950  => x"f3", 951  => x"00", 952  => x"86", 953  => x"00", 954  => x"7c", 955  => x"b8", 956  => x"c3", 957  => x"01", 958  => x"00", 959  => x"00",
      960  => x"88", 961  => x"00", 962  => x"00", 963  => x"00", 964  => x"00", 965  => x"00", 966  => x"00", 967  => x"00", 968  => x"80", 969  => x"00", 970  => x"04", 971  => x"00", 972  => x"00", 973  => x"00", 974  => x"00", 975  => x"00",
      976  => x"70", 977  => x"00", 978  => x"00", 979  => x"00", 980  => x"00", 981  => x"00", 982  => x"00", 983  => x"00", 984  => x"60", 985  => x"00", 986  => x"04", 987  => x"00", 988  => x"00", 989  => x"00", 990  => x"00", 991  => x"00",
      992  => x"00", 993  => x"00", 994  => x"00", 995  => x"00", 996  => x"00", 997  => x"00", 998  => x"00", 999  => x"00", 1000 => x"00", 1001 => x"00", 1002 => x"00", 1003 => x"00", 1004 => x"00", 1005 => x"00", 1006 => x"00", 1007 => x"00",
      1008 => x"00", 1009 => x"00", 1010 => x"00", 1011 => x"00", 1012 => x"00", 1013 => x"00", 1014 => x"00", 1015 => x"00", 1016 => x"00", 1017 => x"00", 1018 => x"00", 1019 => x"00", 1020 => x"00", 1021 => x"00", 1022 => x"00", 1023 => x"00",
      --init code
      1024 => x"ae",
      1025 => x"d5",
      1026 => x"80",
      1027 => x"a8",
      1028 => x"3f",
      1029 => x"d3",
      1030 => x"00",
      1031 => x"40",
      1032 => x"8d",
      1033 => x"14",
      1034 => x"20",
      1035 => x"00",
      1036 => x"a1",
      1037 => x"c8",
      1038 => x"da",
      1039 => x"12",
      1040 => x"81",
      1041 => x"cf",
      1042 => x"d9",
      1043 => x"f1",
      1044 => x"db",
      1045 => x"40",
      1046 => x"a4",
      1047 => x"a6",
      1048 => x"af",
      1049 => x"21",
      1050 => x"00",
      1051 => x"7f",
      1052 => x"22",
      1053 => x"00",
      1054 => x"07",
      others	=> x"00"
   );
   signal program : array_type;
   signal const0 : std_logic := '0';
begin
   
   process(const0)
   begin
      for i in 0 to 1023 loop
         program(i*2) <= prog_instr(i)(15 downto 8);
         program(i*2 + 1) <= prog_instr(i)(7 downto 0);
      end loop;
      for i in 0 to 2047 loop
         program(i + 2048) <= prog_data(i);
      end loop;
   end process;
   data_out <= program(to_integer(unsigned(addr)));
   out_ctl <= '1' when (sel = '1') else '0';

end behavioral;

